`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    18:36:42 03/19/2014 
// Design Name: 
// Module Name:    Memory 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Memory(
				input push,
				input [31:0] addr,
				input WR,
				input IR_DR,
				input [31:0] MDataIn,
				input clk,
				input reset,
				output [31:0] IR,
				output [31:0] DR,
				output [7:0] outans,
				output [3:0] outnumber,
				output [31:0] inter_addr
    );

	reg [31:0] code [18:0];
	reg [31:0] data [7:0];
	
	reg rstuse =1;
	
	reg [31:0] i =0;
	reg [31:0] d =0;
	
	reg [2:0] count =0;
	reg [7:0] aout =0;
	
	assign outans = aout;
	assign outnumber =count;
	assign inter_addr = 11;		//�ж�������ͷ
	
	always @(posedge push)
	begin
		count =count+1;
	end

	
	always @(posedge push)
	begin
		case(count)
		3'b000:aout = data[1];
		3'b001:aout = data[2];
		3'b010:aout = data[3];
		3'b011:aout = data[4];
		3'b100:aout = data[5];
		3'b101:aout = data[6];
		3'b110:aout = data[7];
		3'b111:aout = data[0];
		endcase
	end
	
	
	always @(posedge clk)
	begin
		if(reset?1:rstuse)
		begin			//   b11111122222333334444455555666666		
		//	code[1] <= 32'b10011100000000000000000000000000;
		//	code[0] <= 32'b00100000001000000000000000000011;
		/*	
			code[0] <= 32'b00000000000000000000000000000000;		//nop
			code[1] <= 32'b00100000010000000000000000000001;		//addi s2,s0,1 
			code[2] <= 32'b00100000001000000000000000000001;		//addi s1,s0,1
			code[3] <= 32'b00010000001000100000000000000001;		//beq  s1,s2,1	
			code[4] <= 32'b00000000011000100000100000100000;		//add  s3,s2,s1
			code[5] <= 32'b00100000011000000000000000001001;		//addi s3,s0,9
			code[6] <= 32'b00000000110000110000100000100000;		//add	 6,3,1
			code[7] <= 32'b00000000110000110001100000100000;		//add	 6,3,3
			code[8] <= 32'b10011100000000000000000000000000;		//halt
			code[9] <= 32'b10011100000000000000000000000000;		//halt

		*/
		/*
			code[0] <= 32'b00000000000000000000000000000000;
			code[1] <= 32'b00100000011000000000000000000101;		//addi s3,s0,5
			code[2] <= 32'b00100000001000000000000000000000;		//addi s1,s0,0
			code[3] <= 32'b00100000101000000000000000000001;		//addi s5,s0,1
			code[4] <= 32'b00000000110000010010100000100000;		//add  s6,s1,s5
			code[5] <= 32'b00000000001001100000000000100000;		//add  s1,s6,s0
			code[6] <= 32'b00000000100000100000100000100000;		//add  s4,s2,s1
			code[7] <= 32'b00000000010001000000000000100000;		//add  s2,s4,s0
			code[8] <= 32'b00010100001000111111111111111011;		//bne  s1,s3,-5
			code[9] <= 32'b10011100000000000000000000000000;		//halt
			code[10] <= 32'b10011100000000000000000000000000;		//halt
		*/

			code[0] <= 32'b00000000000000000000000000000000;		//nop
			code[1] <= 32'b10001100001000000000000000000011;		//lw s1,s0,3
			code[2] <= 32'b10001100010000000000000000000010;		//lw s2,s0,2
			code[3] <= 32'b00000000011000100000100000100000;		//add s3,s2,s1
			code[4] <= 32'b01100000000000000000000000000000;		//interrupt
			code[5] <= 32'b10001100100000000000000000000001;		//lw s4,s0,1
			code[6] <= 32'b00000000101001000001100000100100;		//and s5,s4,s3
			code[7] <= 32'b10101100101000000000000000000000;		//sw s5,s0,0
			code[8] <= 32'b10011100000000000000000000000000;		//halt
			code[9] <= 32'b10011100000000000000000000000000;		//halt
			code[10] <= 32'b10011100000000000000000000000000;		//halt
			code[11] <= 32'b00100000111000000000000010101100;		//addi s7,0xac
			code[12] <= 32'b01101100000000000000000000000000;		//ret

	/*		
			code[0] <= 32'b00000000000000000000000000000000;		//nop
	//		code[1] <= 32'b00100000001000000111111111111111;		//addi s1,s0,2^15-1
			code[1] <= 32'b00100000001000001111111111111111;
	//		code[2] <= 32'b00100000011000000111111111111111;		//addi s2,s0,2^15-1
			code[2] <= 32'b00100000011000001111111111111111;
			code[3] <= 32'b00000000011000100000100000100000;		//add s3,s2,s1
			code[4] <= 32'b00000000010000110000100000100000;		//add s2,s3,s1	
			code[5] <= 32'b00011100000000000000000000000001;		//jo +1
			code[6] <= 32'b00001011111111111111111111111101;		//jmp -3
			code[7] <= 32'b10001100100000000000000000000011;		//lw
			code[8] <= 32'b10101100101000000000000000000000;		//sw s5,s0,0
			code[9] <= 32'b10011100000000000000000000000000;		//halt
			code[10] <= 32'b10011100000000000000000000000000;		//halt
			code[11] <= 32'b00100000111000000000000010101100;		//addi s7,0xac
			code[12] <= 32'b01101100000000000000000000000000;		//ret
*/
			
			
			data[0] <= 32'b00000000000000000000000000000111;		//7
			data[1] <= 32'b00000000000000000000000000001000;		//8
			data[2] <= 32'b00000000000000000000000000001100;		//c
			data[3] <= 32'b00000000000000000000000010101100;		//ac
			data[4] <= 32'b00000000000000000000000000000010;		//2
			data[5] <= 32'b00000000000000000000000000000011;		//3
			data[6] <= 32'b00000000000000000000000000001100;		//c
			data[7] <= 32'b00000000000000000000000000000110;		//6

			
			i <= 32'b00000000000000000000000000000000;
			d <= 32'b00000000000000000000000000000000;
			rstuse<=0;
		end
 
		begin
			case(WR)
			1'b0:		 			//write in
				data[addr] <= MDataIn;
			1'b1:					//read out
				case(IR_DR)
					1'b0:
					begin
					if(addr)
						i <= code[addr];
					else
						i <= code[0];
					end
					1'b1:
					begin
					if(addr)
						d <= data[addr];
					else
						d <= data[0];
					end
				endcase
			endcase
		end
		
	end
	
	assign IR = i;
	assign DR = d;
	

endmodule
